library ieee;
use ieee.std_logic_1164.all;

entity shift1_4_tb is
end entity shift1_4_tb;

architecture bhv of shift1_4_tb is

	constant T_CLK 		: time := 10 ns;
	constant T_RESET 	: time := 25 ns;
	signal	clk_tb		  

begin
	
end architecture bhv;